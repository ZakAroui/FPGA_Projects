library ieee;
use ieee.std_logic_1164.all;
entity decoder is
port (x:in std_logic_vector (3 downto 0);
      y: out std_logic_vector (6 downto 0));
end decoder ;
architecture case_when of decoder is
begin 
 process (x)
 begin 
   case x is 
  when "0000" => y<="1000000";
  when "0001" => y<="1111001";
  when "0010" => y<="0100100";
  when "0011" => y<="0110000";
  when "0100" => y<="0011001";
  when "0101" => y<="0010010";
  when "0110" => y<="0000010";
  when "0111" => y<="1111000";
  when "1000" => y<="0000000";
  when "1001" => y<="0010000";
  when "1010" => y<="0001000";
  when "1011" => y<="0000011";
  when "1100" => y<="1000110";
  when "1101" => y<="0100001";
  when "1110" => y<="0000110";
  when others => y<="0001110";
 end case;
 end process;
end case_when;